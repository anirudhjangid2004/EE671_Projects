magic
tech sky130A
timestamp 1726400728
<< error_p >>
rect 685 100 730 113
<< nmos >>
rect 0 135 15 260
rect 140 135 155 260
rect 280 135 295 260
rect 420 135 435 260
rect 560 135 575 260
rect 700 135 715 260
rect 840 135 855 260
rect 980 135 995 260
rect 1120 135 1135 260
rect 1260 135 1275 260
rect 1400 135 1415 260
rect 0 15 15 57
rect 140 15 155 57
rect 280 15 295 57
rect 420 15 435 57
rect 560 15 575 57
rect 700 15 715 57
rect 840 15 855 57
rect 980 15 995 57
rect 1120 15 1135 57
rect 1260 15 1275 57
rect 1400 15 1415 57
<< ndiff >>
rect -45 245 0 260
rect -45 225 -35 245
rect -10 225 0 245
rect -45 205 0 225
rect -45 185 -35 205
rect -10 185 0 205
rect -45 165 0 185
rect -45 145 -35 165
rect -10 145 0 165
rect -45 135 0 145
rect 15 245 60 260
rect 15 225 25 245
rect 50 225 60 245
rect 15 205 60 225
rect 15 185 25 205
rect 50 185 60 205
rect 15 165 60 185
rect 15 145 25 165
rect 50 145 60 165
rect 15 135 60 145
rect 95 245 140 260
rect 95 225 105 245
rect 130 225 140 245
rect 95 205 140 225
rect 95 185 105 205
rect 130 185 140 205
rect 95 165 140 185
rect 95 145 105 165
rect 130 145 140 165
rect 95 135 140 145
rect 155 245 200 260
rect 155 225 165 245
rect 190 225 200 245
rect 155 205 200 225
rect 155 185 165 205
rect 190 185 200 205
rect 155 165 200 185
rect 155 145 165 165
rect 190 145 200 165
rect 155 135 200 145
rect 235 245 280 260
rect 235 225 245 245
rect 270 225 280 245
rect 235 205 280 225
rect 235 185 245 205
rect 270 185 280 205
rect 235 165 280 185
rect 235 145 245 165
rect 270 145 280 165
rect 235 135 280 145
rect 295 245 340 260
rect 295 225 305 245
rect 330 225 340 245
rect 295 205 340 225
rect 295 185 305 205
rect 330 185 340 205
rect 295 165 340 185
rect 295 145 305 165
rect 330 145 340 165
rect 295 135 340 145
rect 375 245 420 260
rect 375 225 385 245
rect 410 225 420 245
rect 375 205 420 225
rect 375 185 385 205
rect 410 185 420 205
rect 375 165 420 185
rect 375 145 385 165
rect 410 145 420 165
rect 375 135 420 145
rect 435 245 480 260
rect 435 225 445 245
rect 470 225 480 245
rect 435 205 480 225
rect 435 185 445 205
rect 470 185 480 205
rect 435 165 480 185
rect 435 145 445 165
rect 470 145 480 165
rect 435 135 480 145
rect 515 245 560 260
rect 515 225 525 245
rect 550 225 560 245
rect 515 205 560 225
rect 515 185 525 205
rect 550 185 560 205
rect 515 165 560 185
rect 515 145 525 165
rect 550 145 560 165
rect 515 135 560 145
rect 575 245 620 260
rect 575 225 585 245
rect 610 225 620 245
rect 575 205 620 225
rect 575 185 585 205
rect 610 185 620 205
rect 575 165 620 185
rect 575 145 585 165
rect 610 145 620 165
rect 575 135 620 145
rect 655 245 700 260
rect 655 225 665 245
rect 690 225 700 245
rect 655 205 700 225
rect 655 185 665 205
rect 690 185 700 205
rect 655 165 700 185
rect 655 145 665 165
rect 690 145 700 165
rect 655 135 700 145
rect 715 245 760 260
rect 715 225 725 245
rect 750 225 760 245
rect 715 205 760 225
rect 715 185 725 205
rect 750 185 760 205
rect 715 165 760 185
rect 715 145 725 165
rect 750 145 760 165
rect 715 135 760 145
rect 795 245 840 260
rect 795 225 805 245
rect 830 225 840 245
rect 795 205 840 225
rect 795 185 805 205
rect 830 185 840 205
rect 795 165 840 185
rect 795 145 805 165
rect 830 145 840 165
rect 795 135 840 145
rect 855 245 900 260
rect 855 225 865 245
rect 890 225 900 245
rect 855 205 900 225
rect 855 185 865 205
rect 890 185 900 205
rect 855 165 900 185
rect 855 145 865 165
rect 890 145 900 165
rect 855 135 900 145
rect 935 245 980 260
rect 935 225 945 245
rect 970 225 980 245
rect 935 205 980 225
rect 935 185 945 205
rect 970 185 980 205
rect 935 165 980 185
rect 935 145 945 165
rect 970 145 980 165
rect 935 135 980 145
rect 995 245 1040 260
rect 995 225 1005 245
rect 1030 225 1040 245
rect 995 205 1040 225
rect 995 185 1005 205
rect 1030 185 1040 205
rect 995 165 1040 185
rect 995 145 1005 165
rect 1030 145 1040 165
rect 995 135 1040 145
rect 1075 245 1120 260
rect 1075 225 1085 245
rect 1110 225 1120 245
rect 1075 205 1120 225
rect 1075 185 1085 205
rect 1110 185 1120 205
rect 1075 165 1120 185
rect 1075 145 1085 165
rect 1110 145 1120 165
rect 1075 135 1120 145
rect 1135 245 1180 260
rect 1135 225 1145 245
rect 1170 225 1180 245
rect 1135 205 1180 225
rect 1135 185 1145 205
rect 1170 185 1180 205
rect 1135 165 1180 185
rect 1135 145 1145 165
rect 1170 145 1180 165
rect 1135 135 1180 145
rect 1215 245 1260 260
rect 1215 225 1225 245
rect 1250 225 1260 245
rect 1215 205 1260 225
rect 1215 185 1225 205
rect 1250 185 1260 205
rect 1215 165 1260 185
rect 1215 145 1225 165
rect 1250 145 1260 165
rect 1215 135 1260 145
rect 1275 245 1320 260
rect 1275 225 1285 245
rect 1310 225 1320 245
rect 1275 205 1320 225
rect 1275 185 1285 205
rect 1310 185 1320 205
rect 1275 165 1320 185
rect 1275 145 1285 165
rect 1310 145 1320 165
rect 1275 135 1320 145
rect 1355 245 1400 260
rect 1355 225 1365 245
rect 1390 225 1400 245
rect 1355 205 1400 225
rect 1355 185 1365 205
rect 1390 185 1400 205
rect 1355 165 1400 185
rect 1355 145 1365 165
rect 1390 145 1400 165
rect 1355 135 1400 145
rect 1415 245 1460 260
rect 1415 225 1425 245
rect 1450 225 1460 245
rect 1415 205 1460 225
rect 1415 185 1425 205
rect 1450 185 1460 205
rect 1415 165 1460 185
rect 1415 145 1425 165
rect 1450 145 1460 165
rect 1415 135 1460 145
rect -45 45 0 57
rect -45 25 -35 45
rect -10 25 0 45
rect -45 15 0 25
rect 15 45 60 57
rect 15 25 25 45
rect 50 25 60 45
rect 15 15 60 25
rect 95 45 140 57
rect 95 25 105 45
rect 130 25 140 45
rect 95 15 140 25
rect 155 45 200 57
rect 155 25 165 45
rect 190 25 200 45
rect 155 15 200 25
rect 235 45 280 57
rect 235 25 245 45
rect 270 25 280 45
rect 235 15 280 25
rect 295 45 340 57
rect 295 25 305 45
rect 330 25 340 45
rect 295 15 340 25
rect 375 45 420 57
rect 375 25 385 45
rect 410 25 420 45
rect 375 15 420 25
rect 435 45 480 57
rect 435 25 445 45
rect 470 25 480 45
rect 435 15 480 25
rect 515 45 560 57
rect 515 25 525 45
rect 550 25 560 45
rect 515 15 560 25
rect 575 45 620 57
rect 575 25 585 45
rect 610 25 620 45
rect 575 15 620 25
rect 655 45 700 57
rect 655 25 665 45
rect 690 25 700 45
rect 655 15 700 25
rect 715 45 760 57
rect 715 25 725 45
rect 750 25 760 45
rect 715 15 760 25
rect 795 45 840 57
rect 795 25 805 45
rect 830 25 840 45
rect 795 15 840 25
rect 855 45 900 57
rect 855 25 865 45
rect 890 25 900 45
rect 855 15 900 25
rect 935 45 980 57
rect 935 25 945 45
rect 970 25 980 45
rect 935 15 980 25
rect 995 45 1040 57
rect 995 25 1005 45
rect 1030 25 1040 45
rect 995 15 1040 25
rect 1075 45 1120 57
rect 1075 25 1085 45
rect 1110 25 1120 45
rect 1075 15 1120 25
rect 1135 45 1180 57
rect 1135 25 1145 45
rect 1170 25 1180 45
rect 1135 15 1180 25
rect 1215 45 1260 57
rect 1215 25 1225 45
rect 1250 25 1260 45
rect 1215 15 1260 25
rect 1275 45 1320 57
rect 1275 25 1285 45
rect 1310 25 1320 45
rect 1275 15 1320 25
rect 1355 45 1400 57
rect 1355 25 1365 45
rect 1390 25 1400 45
rect 1355 15 1400 25
rect 1415 45 1460 57
rect 1415 25 1425 45
rect 1450 25 1460 45
rect 1415 15 1460 25
<< ndiffc >>
rect -35 225 -10 245
rect -35 185 -10 205
rect -35 145 -10 165
rect 25 225 50 245
rect 25 185 50 205
rect 25 145 50 165
rect 105 225 130 245
rect 105 185 130 205
rect 105 145 130 165
rect 165 225 190 245
rect 165 185 190 205
rect 165 145 190 165
rect 245 225 270 245
rect 245 185 270 205
rect 245 145 270 165
rect 305 225 330 245
rect 305 185 330 205
rect 305 145 330 165
rect 385 225 410 245
rect 385 185 410 205
rect 385 145 410 165
rect 445 225 470 245
rect 445 185 470 205
rect 445 145 470 165
rect 525 225 550 245
rect 525 185 550 205
rect 525 145 550 165
rect 585 225 610 245
rect 585 185 610 205
rect 585 145 610 165
rect 665 225 690 245
rect 665 185 690 205
rect 665 145 690 165
rect 725 225 750 245
rect 725 185 750 205
rect 725 145 750 165
rect 805 225 830 245
rect 805 185 830 205
rect 805 145 830 165
rect 865 225 890 245
rect 865 185 890 205
rect 865 145 890 165
rect 945 225 970 245
rect 945 185 970 205
rect 945 145 970 165
rect 1005 225 1030 245
rect 1005 185 1030 205
rect 1005 145 1030 165
rect 1085 225 1110 245
rect 1085 185 1110 205
rect 1085 145 1110 165
rect 1145 225 1170 245
rect 1145 185 1170 205
rect 1145 145 1170 165
rect 1225 225 1250 245
rect 1225 185 1250 205
rect 1225 145 1250 165
rect 1285 225 1310 245
rect 1285 185 1310 205
rect 1285 145 1310 165
rect 1365 225 1390 245
rect 1365 185 1390 205
rect 1365 145 1390 165
rect 1425 225 1450 245
rect 1425 185 1450 205
rect 1425 145 1450 165
rect -35 25 -10 45
rect 25 25 50 45
rect 105 25 130 45
rect 165 25 190 45
rect 245 25 270 45
rect 305 25 330 45
rect 385 25 410 45
rect 445 25 470 45
rect 525 25 550 45
rect 585 25 610 45
rect 665 25 690 45
rect 725 25 750 45
rect 805 25 830 45
rect 865 25 890 45
rect 945 25 970 45
rect 1005 25 1030 45
rect 1085 25 1110 45
rect 1145 25 1170 45
rect 1225 25 1250 45
rect 1285 25 1310 45
rect 1365 25 1390 45
rect 1425 25 1450 45
<< psubdiff >>
rect -100 245 -45 260
rect -100 225 -85 245
rect -60 225 -45 245
rect -100 205 -45 225
rect -100 185 -85 205
rect -60 185 -45 205
rect -100 165 -45 185
rect -100 145 -85 165
rect -60 145 -45 165
rect -100 135 -45 145
rect -100 45 -45 57
rect -100 25 -85 45
rect -60 25 -45 45
rect -100 15 -45 25
<< psubdiffcont >>
rect -85 225 -60 245
rect -85 185 -60 205
rect -85 145 -60 165
rect -85 25 -60 45
<< poly >>
rect 0 260 15 273
rect 140 260 155 273
rect 280 260 295 273
rect 420 260 435 273
rect 560 260 575 273
rect 700 260 715 273
rect 840 260 855 273
rect 980 260 995 273
rect 1120 260 1135 273
rect 1260 260 1275 273
rect 1400 260 1415 273
rect 0 57 15 135
rect 140 120 155 135
rect 280 110 295 135
rect 420 110 435 135
rect 560 120 575 135
rect 700 125 715 135
rect 255 104 295 110
rect 255 87 265 104
rect 286 87 295 104
rect 255 80 295 87
rect 395 104 435 110
rect 395 87 405 104
rect 426 87 435 104
rect 685 100 730 125
rect 840 110 855 135
rect 980 110 995 135
rect 815 104 855 110
rect 395 80 435 87
rect 140 57 155 70
rect 280 57 295 80
rect 420 57 435 80
rect 560 57 575 70
rect 685 67 730 92
rect 815 87 825 104
rect 846 87 855 104
rect 815 80 855 87
rect 955 104 995 110
rect 1120 127 1135 135
rect 1120 108 1195 127
rect 955 87 965 104
rect 986 87 995 104
rect 1156 97 1195 108
rect 955 80 995 87
rect 700 57 715 67
rect 840 57 855 80
rect 980 57 995 80
rect 1060 85 1099 95
rect 1060 66 1135 85
rect 1120 57 1135 66
rect 1260 57 1275 135
rect 1400 110 1415 135
rect 1375 103 1415 110
rect 1375 86 1385 103
rect 1406 86 1415 103
rect 1375 80 1415 86
rect 1400 57 1415 80
rect 0 0 15 15
rect 140 0 155 15
rect 280 0 295 15
rect 420 0 435 15
rect 560 0 575 15
rect 700 0 715 15
rect 840 0 855 15
rect 980 0 995 15
rect 1120 0 1135 15
rect 1260 0 1275 15
rect 1400 0 1415 15
<< polycont >>
rect 265 87 286 104
rect 405 87 426 104
rect 825 87 846 104
rect 965 87 986 104
rect 1385 86 1406 103
<< locali >>
rect -100 280 1460 300
rect -90 245 -57 280
rect -90 225 -85 245
rect -60 225 -57 245
rect -90 205 -57 225
rect -90 185 -85 205
rect -60 185 -57 205
rect -90 165 -57 185
rect -90 145 -85 165
rect -60 145 -57 165
rect -90 135 -57 145
rect -40 245 -5 280
rect -40 225 -35 245
rect -10 225 -5 245
rect -40 205 -5 225
rect -40 185 -35 205
rect -10 185 -5 205
rect -40 165 -5 185
rect -40 145 -35 165
rect -10 145 -5 165
rect -40 135 -5 145
rect 20 245 55 260
rect 100 245 135 260
rect 20 225 25 245
rect 50 225 105 245
rect 130 225 135 245
rect 20 205 55 225
rect 100 205 135 225
rect 20 185 25 205
rect 50 185 105 205
rect 130 185 135 205
rect 20 165 55 185
rect 100 165 135 185
rect 20 145 25 165
rect 50 145 105 165
rect 130 145 135 165
rect 20 135 55 145
rect 100 135 135 145
rect 160 245 195 260
rect 160 225 165 245
rect 190 225 195 245
rect 160 205 195 225
rect 160 185 165 205
rect 190 185 195 205
rect 160 165 195 185
rect 160 145 165 165
rect 190 145 195 165
rect 160 135 195 145
rect 240 245 275 280
rect 240 225 245 245
rect 270 225 275 245
rect 240 205 275 225
rect 240 185 245 205
rect 270 185 275 205
rect 240 165 275 185
rect 240 145 245 165
rect 270 145 275 165
rect 240 135 275 145
rect 300 245 335 260
rect 300 225 305 245
rect 330 225 335 245
rect 300 205 335 225
rect 300 185 305 205
rect 330 185 335 205
rect 300 165 335 185
rect 300 145 305 165
rect 330 145 335 165
rect 300 135 335 145
rect 380 245 415 280
rect 380 225 385 245
rect 410 225 415 245
rect 380 205 415 225
rect 380 185 385 205
rect 410 185 415 205
rect 380 165 415 185
rect 380 145 385 165
rect 410 145 415 165
rect 380 135 415 145
rect 440 245 475 260
rect 520 245 555 260
rect 440 225 445 245
rect 470 225 525 245
rect 550 225 555 245
rect 440 205 475 225
rect 520 205 555 225
rect 440 185 445 205
rect 470 185 525 205
rect 550 185 555 205
rect 440 165 475 185
rect 520 165 555 185
rect 440 145 445 165
rect 470 145 525 165
rect 550 145 555 165
rect 440 135 475 145
rect 520 135 555 145
rect 580 245 615 260
rect 580 225 585 245
rect 610 225 615 245
rect 580 205 615 225
rect 580 185 585 205
rect 610 185 615 205
rect 580 165 615 185
rect 580 145 585 165
rect 610 145 615 165
rect 580 135 615 145
rect 660 245 695 260
rect 660 225 665 245
rect 690 225 695 245
rect 660 205 695 225
rect 660 185 665 205
rect 690 185 695 205
rect 660 165 695 185
rect 660 145 665 165
rect 690 145 695 165
rect 660 135 695 145
rect 720 245 755 260
rect 720 225 725 245
rect 750 225 755 245
rect 720 205 755 225
rect 720 185 725 205
rect 750 185 755 205
rect 720 165 755 185
rect 720 145 725 165
rect 750 145 755 165
rect 720 135 755 145
rect 800 245 835 280
rect 800 225 805 245
rect 830 225 835 245
rect 800 205 835 225
rect 800 185 805 205
rect 830 185 835 205
rect 800 165 835 185
rect 800 145 805 165
rect 830 145 835 165
rect 800 135 835 145
rect 860 245 895 260
rect 860 225 865 245
rect 890 225 895 245
rect 860 205 895 225
rect 860 185 865 205
rect 890 185 895 205
rect 860 165 895 185
rect 860 145 865 165
rect 890 145 895 165
rect 860 135 895 145
rect 940 245 975 280
rect 940 225 945 245
rect 970 225 975 245
rect 940 205 975 225
rect 940 185 945 205
rect 970 185 975 205
rect 940 165 975 185
rect 940 145 945 165
rect 970 145 975 165
rect 940 135 975 145
rect 1000 245 1035 260
rect 1080 245 1115 260
rect 1000 225 1005 245
rect 1030 225 1085 245
rect 1110 225 1115 245
rect 1000 205 1035 225
rect 1080 205 1115 225
rect 1000 185 1005 205
rect 1030 185 1085 205
rect 1110 185 1115 205
rect 1000 165 1035 185
rect 1080 165 1115 185
rect 1000 145 1005 165
rect 1030 145 1085 165
rect 1110 145 1115 165
rect 1000 135 1035 145
rect 1080 135 1115 145
rect 1140 245 1175 260
rect 1140 225 1145 245
rect 1170 225 1175 245
rect 1140 205 1175 225
rect 1140 185 1145 205
rect 1170 185 1175 205
rect 1140 165 1175 185
rect 1140 145 1145 165
rect 1170 145 1175 165
rect 1140 137 1175 145
rect 1220 245 1255 280
rect 1220 225 1225 245
rect 1250 225 1255 245
rect 1220 205 1255 225
rect 1220 185 1225 205
rect 1250 185 1255 205
rect 1220 165 1255 185
rect 1220 145 1225 165
rect 1250 145 1255 165
rect 1220 135 1255 145
rect 1280 245 1315 260
rect 1280 225 1285 245
rect 1310 225 1315 245
rect 1280 205 1315 225
rect 1280 185 1285 205
rect 1310 185 1315 205
rect 1280 165 1315 185
rect 1280 145 1285 165
rect 1310 145 1315 165
rect 1280 135 1315 145
rect 1360 245 1395 280
rect 1360 225 1365 245
rect 1390 225 1395 245
rect 1360 205 1395 225
rect 1360 185 1365 205
rect 1390 185 1395 205
rect 1360 165 1395 185
rect 1360 145 1365 165
rect 1390 145 1395 165
rect 1360 135 1395 145
rect 1420 245 1455 260
rect 1420 225 1425 245
rect 1450 225 1455 245
rect 1420 205 1455 225
rect 1420 185 1425 205
rect 1450 185 1455 205
rect 1420 165 1455 185
rect 1420 145 1425 165
rect 1450 145 1455 165
rect 1420 135 1455 145
rect 35 57 55 135
rect 175 105 195 135
rect 255 105 295 110
rect 175 104 295 105
rect 175 87 265 104
rect 286 87 295 104
rect 175 85 295 87
rect 175 57 195 85
rect 255 80 295 85
rect 315 105 335 135
rect 395 105 435 110
rect 315 104 435 105
rect 315 87 405 104
rect 426 87 435 104
rect 315 85 435 87
rect 315 57 335 85
rect 395 80 435 85
rect 455 57 475 135
rect 660 57 680 135
rect 735 105 755 135
rect 815 105 855 110
rect 735 104 855 105
rect 735 87 825 104
rect 846 87 855 104
rect 735 85 855 87
rect 735 57 755 85
rect 815 80 855 85
rect 875 105 895 135
rect 955 105 995 110
rect 875 104 995 105
rect 875 87 965 104
rect 986 87 995 104
rect 875 85 995 87
rect -90 45 -57 57
rect -90 25 -85 45
rect -60 25 -57 45
rect -90 -5 -57 25
rect -40 45 -5 57
rect -40 25 -35 45
rect -10 25 -5 45
rect -40 -5 -5 25
rect 20 45 55 57
rect 100 45 135 57
rect 20 25 25 45
rect 50 25 105 45
rect 130 25 135 45
rect 20 15 55 25
rect 100 15 135 25
rect 160 45 195 57
rect 160 25 165 45
rect 190 25 195 45
rect 160 15 195 25
rect 240 45 275 57
rect 240 25 245 45
rect 270 25 275 45
rect 240 -5 275 25
rect 300 45 335 57
rect 300 25 305 45
rect 330 25 335 45
rect 300 15 335 25
rect 380 45 415 57
rect 380 25 385 45
rect 410 25 415 45
rect 380 -5 415 25
rect 440 45 475 57
rect 520 45 555 57
rect 440 25 445 45
rect 470 25 525 45
rect 550 25 555 45
rect 440 15 475 25
rect 520 15 555 25
rect 580 45 615 57
rect 580 25 585 45
rect 610 25 615 45
rect 580 15 615 25
rect 660 45 695 57
rect 660 25 665 45
rect 690 25 695 45
rect 660 15 695 25
rect 720 45 755 57
rect 875 55 895 85
rect 955 80 995 85
rect 1015 55 1035 135
rect 1160 117 1190 120
rect 1160 100 1165 117
rect 1185 100 1190 117
rect 1160 97 1190 100
rect 1065 92 1095 95
rect 1065 75 1070 92
rect 1090 75 1095 92
rect 1065 73 1095 75
rect 1295 57 1315 135
rect 1375 103 1415 110
rect 1375 86 1385 103
rect 1406 86 1415 103
rect 1375 80 1415 86
rect 1435 105 1455 135
rect 1435 85 1475 105
rect 1435 57 1455 85
rect 720 25 725 45
rect 750 25 755 45
rect 720 15 755 25
rect 800 45 835 55
rect 800 25 805 45
rect 830 25 835 45
rect 800 -5 835 25
rect 860 45 895 55
rect 860 25 865 45
rect 890 25 895 45
rect 860 15 895 25
rect 940 45 975 55
rect 940 25 945 45
rect 970 25 975 45
rect 940 -5 975 25
rect 1000 45 1035 55
rect 1080 45 1115 55
rect 1000 25 1005 45
rect 1030 25 1085 45
rect 1110 25 1115 45
rect 1000 15 1035 25
rect 1080 15 1115 25
rect 1140 45 1175 57
rect 1140 25 1145 45
rect 1170 25 1175 45
rect 1140 15 1175 25
rect 1220 45 1255 57
rect 1220 25 1225 45
rect 1250 25 1255 45
rect 1220 -5 1255 25
rect 1280 45 1315 57
rect 1280 25 1285 45
rect 1310 25 1315 45
rect 1280 15 1315 25
rect 1360 45 1395 57
rect 1360 25 1365 45
rect 1390 25 1395 45
rect 1360 -5 1395 25
rect 1420 45 1455 57
rect 1420 25 1425 45
rect 1450 25 1455 45
rect 1420 15 1455 25
rect -100 -25 1460 -5
<< viali >>
rect 165 225 190 245
rect 305 145 330 165
rect 585 225 610 245
rect 665 145 690 165
rect 725 225 750 245
rect 1005 145 1030 165
rect 1145 225 1170 245
rect 165 25 190 45
rect 585 25 610 45
rect 1165 100 1185 117
rect 1070 75 1090 92
rect 1385 86 1406 103
rect 725 25 750 45
rect 1145 25 1170 45
<< metal1 >>
rect 160 245 615 255
rect 160 225 165 245
rect 190 225 585 245
rect 610 225 615 245
rect 160 215 615 225
rect 720 245 1175 255
rect 720 225 725 245
rect 750 225 1145 245
rect 1170 225 1175 245
rect 720 215 1175 225
rect 300 165 695 175
rect 300 145 305 165
rect 330 145 665 165
rect 690 145 695 165
rect 300 135 695 145
rect 1000 165 1416 175
rect 1000 145 1005 165
rect 1030 145 1416 165
rect 1000 140 1416 145
rect 1000 139 1100 140
rect 1000 135 1035 139
rect 1215 135 1416 140
rect 1060 117 1200 125
rect 1060 110 1165 117
rect 1156 100 1165 110
rect 1185 110 1200 117
rect 1185 100 1199 110
rect 1156 97 1199 100
rect 1375 103 1416 135
rect 1060 92 1105 95
rect 1060 75 1070 92
rect 1090 80 1105 92
rect 1375 86 1385 103
rect 1406 86 1416 103
rect 1375 80 1416 86
rect 1090 75 1240 80
rect 1060 65 1240 75
rect 160 45 615 55
rect 160 25 165 45
rect 190 25 585 45
rect 610 25 615 45
rect 160 15 615 25
rect 720 45 1175 51
rect 720 25 725 45
rect 750 25 1145 45
rect 1170 25 1175 45
rect 720 15 1175 25
<< end >>
