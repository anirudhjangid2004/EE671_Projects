magic
tech sky130A
timestamp 1726353994
<< error_p >>
rect -80 57 -68 59
rect -92 35 -90 47
<< nwell >>
rect -110 281 -25 359
rect -110 117 920 281
<< nmos >>
rect 0 15 15 57
rect 140 15 155 57
rect 280 15 295 57
rect 420 15 435 57
rect 560 15 575 57
rect 700 15 715 57
rect 840 15 855 57
<< pmos >>
rect 0 135 15 260
rect 140 135 155 260
rect 280 135 295 260
rect 420 135 435 260
rect 560 135 575 260
rect 700 135 715 260
rect 840 135 855 260
<< ndiff >>
rect -45 45 0 57
rect -45 25 -35 45
rect -10 25 0 45
rect -45 15 0 25
rect 15 45 60 57
rect 15 25 25 45
rect 50 25 60 45
rect 15 15 60 25
rect 95 45 140 57
rect 95 25 105 45
rect 130 25 140 45
rect 95 15 140 25
rect 155 45 200 57
rect 155 25 165 45
rect 190 25 200 45
rect 155 15 200 25
rect 235 45 280 57
rect 235 25 245 45
rect 270 25 280 45
rect 235 15 280 25
rect 295 45 340 57
rect 295 25 305 45
rect 330 25 340 45
rect 295 15 340 25
rect 375 45 420 57
rect 375 25 385 45
rect 410 25 420 45
rect 375 15 420 25
rect 435 45 480 57
rect 435 25 445 45
rect 470 25 480 45
rect 435 15 480 25
rect 515 45 560 57
rect 515 25 525 45
rect 550 25 560 45
rect 515 15 560 25
rect 575 45 620 57
rect 575 25 585 45
rect 610 25 620 45
rect 575 15 620 25
rect 655 45 700 57
rect 655 25 665 45
rect 690 25 700 45
rect 655 15 700 25
rect 715 45 760 57
rect 715 25 725 45
rect 750 25 760 45
rect 715 15 760 25
rect 795 45 840 57
rect 795 25 805 45
rect 830 25 840 45
rect 795 15 840 25
rect 855 45 900 57
rect 855 25 865 45
rect 890 25 900 45
rect 855 15 900 25
<< pdiff >>
rect -45 245 0 260
rect -45 225 -35 245
rect -10 225 0 245
rect -45 205 0 225
rect -45 185 -35 205
rect -10 185 0 205
rect -45 165 0 185
rect -45 145 -35 165
rect -10 145 0 165
rect -45 135 0 145
rect 15 245 60 260
rect 15 225 25 245
rect 50 225 60 245
rect 15 205 60 225
rect 15 185 25 205
rect 50 185 60 205
rect 15 165 60 185
rect 15 145 25 165
rect 50 145 60 165
rect 15 135 60 145
rect 95 245 140 260
rect 95 225 105 245
rect 130 225 140 245
rect 95 205 140 225
rect 95 185 105 205
rect 130 185 140 205
rect 95 165 140 185
rect 95 145 105 165
rect 130 145 140 165
rect 95 135 140 145
rect 155 245 200 260
rect 155 225 165 245
rect 190 225 200 245
rect 155 205 200 225
rect 155 185 165 205
rect 190 185 200 205
rect 155 165 200 185
rect 155 145 165 165
rect 190 145 200 165
rect 155 135 200 145
rect 235 245 280 260
rect 235 225 245 245
rect 270 225 280 245
rect 235 205 280 225
rect 235 185 245 205
rect 270 185 280 205
rect 235 165 280 185
rect 235 145 245 165
rect 270 145 280 165
rect 235 135 280 145
rect 295 245 340 260
rect 295 225 305 245
rect 330 225 340 245
rect 295 205 340 225
rect 295 185 305 205
rect 330 185 340 205
rect 295 165 340 185
rect 295 145 305 165
rect 330 145 340 165
rect 295 135 340 145
rect 375 245 420 260
rect 375 225 385 245
rect 410 225 420 245
rect 375 205 420 225
rect 375 185 385 205
rect 410 185 420 205
rect 375 165 420 185
rect 375 145 385 165
rect 410 145 420 165
rect 375 135 420 145
rect 435 245 480 260
rect 435 225 445 245
rect 470 225 480 245
rect 435 205 480 225
rect 435 185 445 205
rect 470 185 480 205
rect 435 165 480 185
rect 435 145 445 165
rect 470 145 480 165
rect 435 135 480 145
rect 515 245 560 260
rect 515 225 525 245
rect 550 225 560 245
rect 515 205 560 225
rect 515 185 525 205
rect 550 185 560 205
rect 515 165 560 185
rect 515 145 525 165
rect 550 145 560 165
rect 515 135 560 145
rect 575 245 620 260
rect 575 225 585 245
rect 610 225 620 245
rect 575 205 620 225
rect 575 185 585 205
rect 610 185 620 205
rect 575 165 620 185
rect 575 145 585 165
rect 610 145 620 165
rect 575 135 620 145
rect 655 245 700 260
rect 655 225 665 245
rect 690 225 700 245
rect 655 205 700 225
rect 655 185 665 205
rect 690 185 700 205
rect 655 165 700 185
rect 655 145 665 165
rect 690 145 700 165
rect 655 135 700 145
rect 715 245 760 260
rect 715 225 725 245
rect 750 225 760 245
rect 715 205 760 225
rect 715 185 725 205
rect 750 185 760 205
rect 715 165 760 185
rect 715 145 725 165
rect 750 145 760 165
rect 715 135 760 145
rect 795 245 840 260
rect 795 225 805 245
rect 830 225 840 245
rect 795 205 840 225
rect 795 185 805 205
rect 830 185 840 205
rect 795 165 840 185
rect 795 145 805 165
rect 830 145 840 165
rect 795 135 840 145
rect 855 245 900 260
rect 855 225 865 245
rect 890 225 900 245
rect 855 205 900 225
rect 855 185 865 205
rect 890 185 900 205
rect 855 165 900 185
rect 855 145 865 165
rect 890 145 900 165
rect 855 135 900 145
<< ndiffc >>
rect -35 25 -10 45
rect 25 25 50 45
rect 105 25 130 45
rect 165 25 190 45
rect 245 25 270 45
rect 305 25 330 45
rect 385 25 410 45
rect 445 25 470 45
rect 525 25 550 45
rect 585 25 610 45
rect 665 25 690 45
rect 725 25 750 45
rect 805 25 830 45
rect 865 25 890 45
<< pdiffc >>
rect -35 225 -10 245
rect -35 185 -10 205
rect -35 145 -10 165
rect 25 225 50 245
rect 25 185 50 205
rect 25 145 50 165
rect 105 225 130 245
rect 105 185 130 205
rect 105 145 130 165
rect 165 225 190 245
rect 165 185 190 205
rect 165 145 190 165
rect 245 225 270 245
rect 245 185 270 205
rect 245 145 270 165
rect 305 225 330 245
rect 305 185 330 205
rect 305 145 330 165
rect 385 225 410 245
rect 385 185 410 205
rect 385 145 410 165
rect 445 225 470 245
rect 445 185 470 205
rect 445 145 470 165
rect 525 225 550 245
rect 525 185 550 205
rect 525 145 550 165
rect 585 225 610 245
rect 585 185 610 205
rect 585 145 610 165
rect 665 225 690 245
rect 665 185 690 205
rect 665 145 690 165
rect 725 225 750 245
rect 725 185 750 205
rect 725 145 750 165
rect 805 225 830 245
rect 805 185 830 205
rect 805 145 830 165
rect 865 225 890 245
rect 865 185 890 205
rect 865 145 890 165
<< psubdiff >>
rect -90 47 -45 57
rect -90 30 -80 47
rect -63 30 -45 47
rect -90 15 -45 30
<< nsubdiff >>
rect -90 135 -45 260
<< psubdiffcont >>
rect -80 30 -63 47
<< poly >>
rect 0 260 15 275
rect 140 260 155 275
rect 280 260 295 275
rect 420 260 435 275
rect 560 260 575 275
rect 700 260 715 275
rect 840 260 855 275
rect 0 80 15 135
rect 140 80 155 135
rect 0 65 155 80
rect 0 57 15 65
rect 140 57 155 65
rect 280 80 295 135
rect 420 80 435 135
rect 280 65 435 80
rect 280 57 295 65
rect 420 57 435 65
rect 560 80 575 135
rect 700 80 715 135
rect 560 65 715 80
rect 560 57 575 65
rect 700 57 715 65
rect 840 57 855 135
rect 0 0 15 15
rect 140 0 155 15
rect 280 0 295 15
rect 420 0 435 15
rect 560 0 575 15
rect 700 0 715 15
rect 840 0 855 15
<< locali >>
rect -90 299 105 300
rect -90 298 -35 299
rect -90 280 -85 298
rect -58 280 -35 298
rect -85 135 -57 280
rect -40 279 -35 280
rect -10 280 105 299
rect 130 280 525 300
rect 550 280 805 300
rect 830 280 905 300
rect -10 279 -5 280
rect -40 245 -5 279
rect -40 225 -35 245
rect -10 225 -5 245
rect -40 205 -5 225
rect -40 185 -35 205
rect -10 185 -5 205
rect -40 165 -5 185
rect -40 145 -35 165
rect -10 145 -5 165
rect -40 135 -5 145
rect 20 245 55 260
rect 20 225 25 245
rect 50 225 55 245
rect 20 205 55 225
rect 20 185 25 205
rect 50 185 55 205
rect 20 165 55 185
rect 20 145 25 165
rect 50 145 55 165
rect 20 115 55 145
rect 100 245 135 280
rect 100 225 105 245
rect 130 225 135 245
rect 100 205 135 225
rect 100 185 105 205
rect 130 185 135 205
rect 100 165 135 185
rect 100 145 105 165
rect 130 145 135 165
rect 100 135 135 145
rect 160 245 195 260
rect 160 225 165 245
rect 190 225 195 245
rect 160 205 195 225
rect 160 185 165 205
rect 190 185 195 205
rect 160 165 195 185
rect 160 145 165 165
rect 190 145 195 165
rect 160 115 195 145
rect 240 245 275 260
rect 240 225 245 245
rect 270 225 275 245
rect 240 205 275 225
rect 240 185 245 205
rect 270 185 275 205
rect 240 165 275 185
rect 240 145 245 165
rect 270 145 275 165
rect 240 115 275 145
rect 300 245 335 260
rect 300 225 305 245
rect 330 225 335 245
rect 300 205 335 225
rect 300 185 305 205
rect 330 185 335 205
rect 300 165 335 185
rect 300 145 305 165
rect 330 145 335 165
rect 300 135 335 145
rect 380 245 415 260
rect 380 225 385 245
rect 410 225 415 245
rect 380 205 415 225
rect 380 185 385 205
rect 410 185 415 205
rect 380 165 415 185
rect 380 145 385 165
rect 410 145 415 165
rect 380 115 415 145
rect 440 245 475 260
rect 440 225 445 245
rect 470 225 475 245
rect 440 205 475 225
rect 440 185 445 205
rect 470 185 475 205
rect 440 165 475 185
rect 440 145 445 165
rect 470 145 475 165
rect 440 135 475 145
rect 520 245 555 280
rect 520 225 525 245
rect 550 225 555 245
rect 520 205 555 225
rect 520 185 525 205
rect 550 185 555 205
rect 520 165 555 185
rect 520 145 525 165
rect 550 145 555 165
rect 520 135 555 145
rect 580 245 615 260
rect 580 225 585 245
rect 610 225 615 245
rect 580 205 615 225
rect 580 185 585 205
rect 610 185 615 205
rect 580 165 615 185
rect 580 145 585 165
rect 610 145 615 165
rect 580 135 615 145
rect 660 245 695 260
rect 660 225 665 245
rect 690 225 695 245
rect 660 205 695 225
rect 660 185 665 205
rect 690 185 695 205
rect 660 165 695 185
rect 660 145 665 165
rect 690 145 695 165
rect 660 135 695 145
rect 720 245 755 260
rect 720 225 725 245
rect 750 225 755 245
rect 720 205 755 225
rect 720 185 725 205
rect 750 185 755 205
rect 720 165 755 185
rect 720 145 725 165
rect 750 145 755 165
rect 720 135 755 145
rect 800 245 835 280
rect 800 225 805 245
rect 830 225 835 245
rect 800 205 835 225
rect 800 185 805 205
rect 830 185 835 205
rect 800 165 835 185
rect 800 145 805 165
rect 830 145 835 165
rect 800 135 835 145
rect 860 245 895 260
rect 860 225 865 245
rect 890 225 895 245
rect 860 205 895 225
rect 860 185 865 205
rect 890 185 895 205
rect 860 165 895 185
rect 860 145 865 165
rect 890 145 895 165
rect 20 95 415 115
rect 520 75 695 95
rect -90 47 -57 57
rect -90 30 -80 47
rect -63 30 -57 47
rect -90 15 -57 30
rect -85 -3 -57 15
rect -85 -23 -84 -3
rect -59 -23 -57 -3
rect -85 -25 -57 -23
rect -40 45 -5 57
rect -40 25 -35 45
rect -10 25 -5 45
rect -40 -5 -5 25
rect 20 45 55 57
rect 20 25 25 45
rect 50 25 55 45
rect 20 15 55 25
rect 100 45 135 57
rect 100 25 105 45
rect 130 25 135 45
rect 100 -5 135 25
rect 160 45 195 57
rect 160 25 165 45
rect 190 25 195 45
rect 160 15 195 25
rect 240 45 275 57
rect 240 25 245 45
rect 270 25 275 45
rect 240 -5 275 25
rect 300 45 335 57
rect 300 25 305 45
rect 330 25 335 45
rect 300 15 335 25
rect 380 45 415 57
rect 380 25 385 45
rect 410 25 415 45
rect 380 -5 415 25
rect 440 45 475 57
rect 440 25 445 45
rect 470 25 475 45
rect 440 15 475 25
rect 520 45 555 75
rect 520 25 525 45
rect 550 25 555 45
rect 520 -5 555 25
rect -40 -25 555 -5
rect 580 45 615 57
rect 580 25 585 45
rect 610 25 615 45
rect 580 -5 615 25
rect 660 45 695 75
rect 660 25 665 45
rect 690 25 695 45
rect 660 15 695 25
rect 720 45 755 57
rect 720 25 725 45
rect 750 25 755 45
rect 720 -5 755 25
rect 800 45 835 55
rect 800 25 805 45
rect 830 25 835 45
rect 800 -5 835 25
rect 860 45 895 145
rect 860 25 865 45
rect 890 25 895 45
rect 860 15 895 25
rect 580 -25 585 -5
rect 610 -25 725 -5
rect 750 -25 805 -5
rect 830 -25 895 -5
<< viali >>
rect -85 280 -58 298
rect -35 279 -10 299
rect 105 280 130 300
rect 525 280 550 300
rect 805 280 830 300
rect 305 225 330 245
rect 305 185 330 205
rect 305 145 330 165
rect 445 225 470 245
rect 445 185 470 205
rect 445 145 470 165
rect 585 225 610 245
rect 585 185 610 205
rect 585 145 610 165
rect -84 -23 -59 -3
rect 25 25 50 45
rect 165 25 190 45
rect 305 25 330 45
rect 445 25 470 45
rect 585 -25 610 -5
rect 725 -25 750 -5
rect 805 -25 830 -5
<< metal1 >>
rect -95 300 910 305
rect -95 299 105 300
rect -95 298 -35 299
rect -95 280 -85 298
rect -58 280 -35 298
rect -95 279 -35 280
rect -10 280 105 299
rect 130 280 525 300
rect 550 280 805 300
rect 830 280 910 300
rect -10 279 910 280
rect -95 275 910 279
rect 300 245 615 260
rect 300 225 305 245
rect 330 225 445 245
rect 470 225 585 245
rect 610 225 615 245
rect 300 205 615 225
rect 300 185 305 205
rect 330 185 445 205
rect 470 185 585 205
rect 610 185 615 205
rect 300 165 615 185
rect 300 145 305 165
rect 330 145 445 165
rect 470 145 585 165
rect 610 145 615 165
rect 300 135 615 145
rect 440 57 475 135
rect 20 45 475 57
rect 20 25 25 45
rect 50 25 165 45
rect 190 25 305 45
rect 330 25 445 45
rect 470 25 475 45
rect 20 15 475 25
rect -95 -3 910 0
rect -95 -23 -84 -3
rect -59 -5 910 -3
rect -59 -23 585 -5
rect -95 -25 585 -23
rect 610 -25 725 -5
rect 750 -25 805 -5
rect 830 -25 910 -5
rect -95 -30 910 -25
<< end >>
