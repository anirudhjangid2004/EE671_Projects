magic
tech sky130A
timestamp 1726353333
<< nwell >>
rect 205 145 810 340
<< nmos >>
rect 325 55 340 105
rect 520 55 535 105
rect 725 55 740 105
<< pmos >>
rect 325 165 340 320
rect 520 165 535 320
rect 725 165 740 320
<< ndiff >>
rect 275 90 325 105
rect 275 70 290 90
rect 310 70 325 90
rect 275 55 325 70
rect 340 90 390 105
rect 340 70 355 90
rect 375 70 390 90
rect 340 55 390 70
rect 470 90 520 105
rect 470 70 487 90
rect 507 70 520 90
rect 470 55 520 70
rect 535 90 585 105
rect 535 70 550 90
rect 570 70 585 90
rect 535 55 585 70
rect 675 90 725 105
rect 675 70 692 90
rect 712 70 725 90
rect 675 55 725 70
rect 740 90 790 105
rect 740 70 755 90
rect 775 70 790 90
rect 740 55 790 70
<< pdiff >>
rect 275 305 325 320
rect 275 180 290 305
rect 310 180 325 305
rect 275 165 325 180
rect 340 305 390 320
rect 340 180 355 305
rect 375 180 390 305
rect 340 165 390 180
rect 470 305 520 320
rect 470 180 485 305
rect 505 180 520 305
rect 470 165 520 180
rect 535 305 585 320
rect 535 180 550 305
rect 570 180 585 305
rect 535 165 585 180
rect 675 305 725 320
rect 675 180 693 305
rect 713 180 725 305
rect 675 165 725 180
rect 740 305 790 320
rect 740 180 755 305
rect 775 180 790 305
rect 740 165 790 180
<< ndiffc >>
rect 290 70 310 90
rect 355 70 375 90
rect 487 70 507 90
rect 550 70 570 90
rect 692 70 712 90
rect 755 70 775 90
<< pdiffc >>
rect 290 180 310 305
rect 355 180 375 305
rect 485 180 505 305
rect 550 180 570 305
rect 693 180 713 305
rect 755 180 775 305
<< psubdiff >>
rect 225 90 275 105
rect 225 70 240 90
rect 260 70 275 90
rect 225 55 275 70
rect 420 90 470 105
rect 420 70 433 90
rect 453 70 470 90
rect 420 55 470 70
rect 625 90 675 105
rect 625 70 638 90
rect 658 70 675 90
rect 625 55 675 70
<< nsubdiff >>
rect 225 305 275 320
rect 225 180 240 305
rect 260 180 275 305
rect 225 165 275 180
rect 420 305 470 320
rect 420 180 435 305
rect 455 180 470 305
rect 420 165 470 180
rect 625 305 675 320
rect 625 180 640 305
rect 660 180 675 305
rect 625 165 675 180
<< psubdiffcont >>
rect 240 70 260 90
rect 433 70 453 90
rect 638 70 658 90
<< nsubdiffcont >>
rect 240 180 260 305
rect 435 180 455 305
rect 640 180 660 305
<< poly >>
rect 325 320 340 335
rect 520 320 535 335
rect 725 320 740 335
rect 325 105 340 165
rect 520 105 535 165
rect 725 105 740 165
rect 325 40 340 55
rect 300 30 340 40
rect 300 10 310 30
rect 330 10 340 30
rect 300 0 340 10
rect 520 5 535 55
rect 725 5 740 55
rect 495 -5 535 5
rect 495 -25 505 -5
rect 525 -25 535 -5
rect 495 -35 535 -25
rect 700 -5 740 5
rect 700 -25 710 -5
rect 730 -25 740 -5
rect 700 -35 740 -25
<< polycont >>
rect 310 10 330 30
rect 505 -25 525 -5
rect 710 -25 730 -5
<< locali >>
rect 560 330 721 350
rect 560 310 580 330
rect 700 310 721 330
rect 230 305 320 310
rect 230 180 240 305
rect 260 180 290 305
rect 310 180 320 305
rect 230 175 320 180
rect 345 305 385 310
rect 345 180 355 305
rect 375 180 385 305
rect 345 175 385 180
rect 425 305 515 310
rect 425 180 435 305
rect 455 180 485 305
rect 505 180 515 305
rect 425 175 515 180
rect 540 305 580 310
rect 540 180 550 305
rect 570 180 580 305
rect 540 175 580 180
rect 630 305 668 310
rect 630 180 640 305
rect 660 180 668 305
rect 630 175 668 180
rect 685 305 721 310
rect 685 180 693 305
rect 713 180 721 305
rect 685 175 721 180
rect 745 305 785 310
rect 745 180 755 305
rect 775 180 785 305
rect 745 175 785 180
rect 365 145 385 175
rect 765 145 785 175
rect 365 125 810 145
rect 560 95 580 125
rect 765 95 785 125
rect 230 90 320 95
rect 230 70 240 90
rect 260 70 290 90
rect 310 70 320 90
rect 230 65 320 70
rect 345 90 385 95
rect 345 70 355 90
rect 375 70 385 90
rect 345 65 385 70
rect 425 90 461 95
rect 425 70 433 90
rect 453 70 461 90
rect 425 65 461 70
rect 479 90 515 95
rect 479 70 487 90
rect 507 70 515 90
rect 479 65 515 70
rect 540 90 580 95
rect 540 70 550 90
rect 570 70 580 90
rect 540 65 580 70
rect 630 90 666 95
rect 630 70 638 90
rect 658 70 666 90
rect 630 65 666 70
rect 684 90 720 95
rect 684 70 692 90
rect 712 70 720 90
rect 684 65 720 70
rect 745 90 785 95
rect 745 70 755 90
rect 775 70 785 90
rect 745 65 785 70
rect 365 45 385 65
rect 495 45 515 65
rect 700 45 720 65
rect 205 30 340 40
rect 205 20 310 30
rect 300 10 310 20
rect 330 10 340 30
rect 365 25 720 45
rect 300 0 340 10
rect 495 -5 535 5
rect 495 -25 505 -5
rect 525 -25 535 -5
rect 495 -35 535 -25
rect 700 -5 740 5
rect 700 -25 710 -5
rect 730 -25 740 -5
rect 700 -35 740 -25
<< viali >>
rect 240 180 260 305
rect 290 180 310 305
rect 435 180 455 305
rect 485 180 505 305
rect 640 180 660 305
rect 240 70 260 90
rect 290 70 310 90
rect 433 70 453 90
rect 638 70 658 90
<< metal1 >>
rect 205 305 810 310
rect 205 180 240 305
rect 260 180 290 305
rect 310 180 435 305
rect 455 180 485 305
rect 505 180 640 305
rect 660 180 810 305
rect 205 175 810 180
rect 205 90 810 95
rect 205 70 240 90
rect 260 70 290 90
rect 310 70 433 90
rect 453 70 638 90
rect 658 70 810 90
rect 205 65 810 70
use inverter  inverter_0
timestamp 1725999080
transform 1 0 120 0 1 55
box -120 -55 85 285
<< labels >>
rlabel metal1 400 243 400 243 7 Vdd
port 3 w
rlabel metal1 605 243 605 243 7 Vdd
port 3 w
rlabel metal1 605 80 605 80 7 Vss
port 2 w
rlabel metal1 400 80 400 80 7 Vss
port 2 w
rlabel metal1 205 80 205 80 7 Vss
port 2 w
rlabel locali 205 29 205 29 7 A
port 1 w
rlabel metal1 205 243 205 243 7 Vdd
port 3 w
<< end >>
